module alu(
    input logic [31:0] source_a, source_b, 
    input logic [1:0] control, 
    output logic [31:0] result, 
    output logic [3:0] flags
    ); 
endmodule
